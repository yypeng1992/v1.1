`timescale 1ns / 1ps
//`include "ddr_define.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    2016/8/4 12:17:58 
// Design Name: 
// Module Name:    ddr_cfg_decoder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ddr_cfg_decoder(
  clk,
  rst_n,
  
  //cfg_network
  cfgid_i,
  cfgfwd_i,
  cfgdata_i,
  cfgreq_i,
  cfgdone_i,
  
  //request info
  request_data_valid_o,     //ȡ�����������Ч��־
  request_pos_1st_o,
  request_pos_2nd_o,
  request_addr_1st_row_o,		//������COP��������
  request_addr_1st_col_o,		//ͬ��..
  request_addr_last_trans_o,//ͬ��..
  
  request_src_type_o,	      //����MCȡָ��    2'b01---256������   2'b10---512������
                            //������ͨȡ����  ������src_a/src_b�ı�ʾ
                            //����copȡָ��   ������src_a/src_b�ı�ʾ
  
  request_cmd_valid_o,			//ȡָ���������Ч��־
  request_cmd_access_addr_o,
  //request_mc_access_addr_o,	//������MCȡ������Ϣ
  //request_cop_access_addr_o,//������COPȡָ��
  

	//cfg info
	cfg_valid_o,
//cfg_get_clu_num_en_o,
//cfg_pos_ok_en_o,
	
	cfg_third_req_o,
	cfg_stream_o,
	cfg_broadcast_o,
	cfg_row_column_o,			//0-��  1-��
	cfg_read_write_o,			//0-��  1-д
	cfg_D2D_flag_o,	
	cfg_ch_cluster_num_o,
	cfg_VR_id_o,					//������������Ĵ������
	cfg_VR_FR_o,
	cfg_ddr_channel_id_o,	//��ַͨ�����
	
	
	//�����cfg info�����ߵ���ʽ�·���32��ddr_channel
  cfg_data_pos0_1st_o,
  cfg_data_pos1_1st_o,
  cfg_data_pos2_1st_o,
  cfg_data_pos3_1st_o,
  cfg_data_pos4_1st_o,
  cfg_data_pos5_1st_o,
  cfg_data_pos6_1st_o,
  cfg_data_pos7_1st_o,
  cfg_data_pos0_2nd_o,
  cfg_data_pos1_2nd_o,
  cfg_data_pos2_2nd_o,
  cfg_data_pos3_2nd_o,
  cfg_data_pos4_2nd_o,
  cfg_data_pos5_2nd_o,
  cfg_data_pos6_2nd_o,
  cfg_data_pos7_2nd_o,
	
  cfg_addr_pos0_1st_o,
  cfg_addr_pos1_1st_o,
  cfg_addr_pos2_1st_o,
  cfg_addr_pos3_1st_o,
  cfg_addr_pos4_1st_o,
  cfg_addr_pos5_1st_o,
  cfg_addr_pos6_1st_o,
  cfg_addr_pos7_1st_o,
  cfg_addr_pos0_2nd_o,
  cfg_addr_pos1_2nd_o,
  cfg_addr_pos2_2nd_o,
  cfg_addr_pos3_2nd_o,
  cfg_addr_pos4_2nd_o,
  cfg_addr_pos5_2nd_o,
  cfg_addr_pos6_2nd_o,
  cfg_addr_pos7_2nd_o,
	
  cfg_start_pos_row_0_o,
  cfg_start_pos_col_0_o,
  cfg_start_pos_row_1_o,
  cfg_start_pos_col_1_o,
  cfg_start_pos_row_2_o,
  cfg_start_pos_col_2_o,
  cfg_start_pos_row_3_o,
  cfg_start_pos_col_3_o,
  cfg_start_pos_row_4_o,
  cfg_start_pos_col_4_o,
  cfg_start_pos_row_5_o,
  cfg_start_pos_col_5_o,
  cfg_start_pos_row_6_o,
  cfg_start_pos_col_6_o,
  cfg_start_pos_row_7_o,
  cfg_start_pos_col_7_o,
	
  cfg_start_addr_o,
  cfg_row_num_1st_o,
  cfg_column_num_1st_o,
  cfg_row_num_2nd_o,
  cfg_column_num_2nd_o,
  cfg_circu_times_o,
  
  /* һ�������������������Ȼ�������,����������ֻ����������,������������ */
	cfg_col_addr_burst_o,	//һ�������м�һ��ַ������Ŀ
	cfg_row_addr_burst_o,	//һ�������м�һ��ַ������Ŀ
	cfg_2nd_addr_burst_o,	//���������м�һ��ַ������Ŀ
	cfg_access_length_burst_o	//���������С--------�涨Ϊ����������е�С���ܸ���
	);
	
	//--------------------------------------------------
	// INPUT && OUTPUT ------- declaration
	//--------------------------------------------------
  input			clk;
  input			rst_n;
  
  //cfg_network
  input			[ 7:0]		cfgid_i;
  input		 		     		cfgfwd_i;
  input			[31:0]		cfgdata_i;
  input		      			cfgreq_i;
  input		      			cfgdone_i;
  
  //request info
  output              request_data_valid_o;
  output    [ 7:0]    request_pos_1st_o;
  output    [ 2:0]    request_pos_2nd_o;
	output    [ 1:0]    request_src_type_o;
  output    [15:0]    request_addr_1st_row_o;
  output    [13:0]    request_addr_1st_col_o;
  output              request_addr_last_trans_o;

	output              request_cmd_valid_o;
	output		[19:0]		request_cmd_access_addr_o;
	//output		[19:0]		request_mc_access_addr_o;
	//output		[11:0]		request_cop_access_addr_o;
	
	
	//cfg info
	output							cfg_valid_o;
//output							cfg_get_clu_num_en_o;
//output							cfg_pos_ok_en_o;
	
	output							cfg_third_req_o;
	output							cfg_stream_o;
	output							cfg_broadcast_o;
	output							cfg_row_column_o;			//0-��  1-��
	output							cfg_read_write_o;			//0-��  1-д
	output							cfg_D2D_flag_o;
	output		[ 2:0]		cfg_ch_cluster_num_o;
	output		[ 8:0]		cfg_VR_id_o;
	output      [ 2:0]      cfg_VR_FR_o;    //// yyp 2016-10-25
	output		[ 4:0]		cfg_ddr_channel_id_o;
	
	
  output		[ 7:0]		cfg_data_pos0_1st_o;
  output		[ 7:0]		cfg_data_pos1_1st_o;
  output		[ 7:0]		cfg_data_pos2_1st_o;
  output		[ 7:0]		cfg_data_pos3_1st_o;
  output		[ 7:0]		cfg_data_pos4_1st_o;
  output		[ 7:0]		cfg_data_pos5_1st_o;
  output		[ 7:0]		cfg_data_pos6_1st_o;
  output		[ 7:0]		cfg_data_pos7_1st_o;
  output		[ 2:0]		cfg_data_pos0_2nd_o;
  output		[ 2:0]		cfg_data_pos1_2nd_o;
  output		[ 2:0]		cfg_data_pos2_2nd_o;
  output		[ 2:0]		cfg_data_pos3_2nd_o;
  output		[ 2:0]		cfg_data_pos4_2nd_o;
  output		[ 2:0]		cfg_data_pos5_2nd_o;
  output		[ 2:0]		cfg_data_pos6_2nd_o;
  output		[ 2:0]		cfg_data_pos7_2nd_o;
	
  output		[ 7:0]		cfg_addr_pos0_1st_o;
  output		[ 7:0]		cfg_addr_pos1_1st_o;
  output		[ 7:0]		cfg_addr_pos2_1st_o;
  output		[ 7:0]		cfg_addr_pos3_1st_o;
  output		[ 7:0]		cfg_addr_pos4_1st_o;
  output		[ 7:0]		cfg_addr_pos5_1st_o;
  output		[ 7:0]		cfg_addr_pos6_1st_o;
  output		[ 7:0]		cfg_addr_pos7_1st_o;
  output		[ 2:0]		cfg_addr_pos0_2nd_o;
  output		[ 2:0]		cfg_addr_pos1_2nd_o;
  output		[ 2:0]		cfg_addr_pos2_2nd_o;
  output		[ 2:0]		cfg_addr_pos3_2nd_o;
  output		[ 2:0]		cfg_addr_pos4_2nd_o;
  output		[ 2:0]		cfg_addr_pos5_2nd_o;
  output		[ 2:0]		cfg_addr_pos6_2nd_o;
  output		[ 2:0]		cfg_addr_pos7_2nd_o;
	
  output	  [15:0]    cfg_start_pos_row_0_o;
  output	  [13:0]    cfg_start_pos_col_0_o;
  output	  [15:0]    cfg_start_pos_row_1_o;
  output	  [13:0]    cfg_start_pos_col_1_o;
  output	  [15:0]    cfg_start_pos_row_2_o;
  output	  [13:0]    cfg_start_pos_col_2_o;
  output	  [15:0]    cfg_start_pos_row_3_o;
  output	  [13:0]    cfg_start_pos_col_3_o;
  output	  [15:0]    cfg_start_pos_row_4_o;
  output	  [13:0]    cfg_start_pos_col_4_o;
  output	  [15:0]    cfg_start_pos_row_5_o;
  output	  [13:0]    cfg_start_pos_col_5_o;
  output	  [15:0]    cfg_start_pos_row_6_o;
  output	  [13:0]    cfg_start_pos_col_6_o;
  output	  [15:0]    cfg_start_pos_row_7_o;
  output	  [13:0]    cfg_start_pos_col_7_o;
	
  output		[29:0]		cfg_start_addr_o;
  output		[15:0]		cfg_row_num_1st_o;
  output		[13:0]		cfg_column_num_1st_o;
  output		[15:0]		cfg_row_num_2nd_o;
  output		[13:0]		cfg_column_num_2nd_o;
  output		[29:0]		cfg_circu_times_o;
	output		[29:0]		cfg_col_addr_burst_o;
	output		[29:0]		cfg_row_addr_burst_o;
	output		[29:0]		cfg_2nd_addr_burst_o;
	output		[29:0]		cfg_access_length_burst_o;
	
	
	//--------------------------------------------------
	// REG && WIRE ------- declaration
	//--------------------------------------------------
	
  //request info
  reg                     request_valid_r;
  reg                     request_cmd_valid_r = 'b0;
  reg		    [ 7:0]    request_pos_1st_r         = 'b0;
  reg		    [ 2:0]    request_pos_2nd_r         = 'b0;
  reg		    [ 1:0]    request_src_type_r        = 'b0;
  reg		    [15:0]    request_addr_1st_row_r    = 'b0;
  reg		    [13:0]    request_addr_1st_col_r    = 'b0;
  reg		              request_addr_last_trans_r = 'b0;
  reg			[19:0]    request_cmd_access_addr_r = 'b0;
  //reg           [19:0]      request_mc_access_addr_r;
	
  
	//cfg info
  reg									cfg_valid_r = 'b0;
//reg									cfg_get_clu_num_en_r;
//reg									cfg_pos_ok_en_r;
  
  reg                 pos_ok_start_pre_r = 'b0; //����cfgid=5
  //reg                 pos_ok_start_en_r;  //����cfgid=6
  
  reg							cfg_third_req_r		= 'b0;
  reg							cfg_stream_r		= 'b0;
  reg							cfg_broadcast_r		= 'b0;
  reg							cfg_row_column_r	= 'b0;
  reg							cfg_read_write_r	= 'b0;
  reg							cfg_D2D_flag_r		= 'b0;
  reg				[ 2:0]		cfg_ch_cluster_num_r= 'b0;
  reg				[ 8:0]		cfg_VR_id_r			= 'b0;
  reg               [ 2:0]      cfg_VR_FR_r			= 'b0;
  reg				[ 4:0]		cfg_ddr_channel_id_r= 'b0;
	
	
  reg				[ 7:0]		cfg_data_pos0_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos1_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos2_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos3_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos4_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos5_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos6_1st_r	= 'b0;
  reg				[ 7:0]		cfg_data_pos7_1st_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos0_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos1_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos2_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos3_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos4_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos5_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos6_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_data_pos7_2nd_r	= 'b0;
	
  reg				[ 7:0]		cfg_addr_pos0_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos1_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos2_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos3_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos4_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos5_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos6_1st_r	= 'b0;
  reg				[ 7:0]		cfg_addr_pos7_1st_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos0_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos1_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos2_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos3_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos4_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos5_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos6_2nd_r	= 'b0;
  reg				[ 2:0]		cfg_addr_pos7_2nd_r	= 'b0;
	
	
  reg				[29:0]		cfg_start_addr_r	= 'b0;
  reg				[15:0]		cfg_row_num_1st_r	= 'b0;
  reg				[13:0]		cfg_column_num_1st_r= 'b0;
  reg				[15:0]		cfg_row_num_2nd_r	= 'b0;
  reg				[13:0]		cfg_column_num_2nd_r= 'b0;
  reg				[29:0]		cfg_circu_times_r	= 'b0;
  reg				[29:0]		cfg_col_addr_burst_r= 'b0;
  reg				[29:0]		cfg_row_addr_burst_r= 'b0;
  reg				[29:0]		cfg_2nd_addr_burst_r= 'b0;
  reg				[29:0]		cfg_access_length_burst_r	= 'b0;
	
	//extra
	reg									cfgreq_r;
	

	//--------------------------------------------------
	// CODE ------- description
	//--------------------------------------------------
	
  //request info ----------------------------
  always@(posedge clk) begin
  	if(!rst_n)
      cfgreq_r <= 1'b0;
    else
      cfgreq_r <= cfgreq_i;
  end
  
  always @(posedge clk) begin
    if(~rst_n)
      request_valid_r <= 1'b0;
    else if(cfgreq_r && cfgdone_i)
      request_valid_r <= 1'b1;
    else
      request_valid_r <= 1'b0;
  end

	//req_0
  always @(posedge clk) begin
    /* if(~rst_n) begin
      request_pos_1st_r  <= 8'b0;
      request_pos_2nd_r  <= 3'b0;
      request_src_type_r <= 2'b0;
    end
    else  */if(cfgreq_i && cfgfwd_i && (cfgid_i == 8'd0)) begin
      request_pos_1st_r  <= cfgdata_i[15: 8];
      request_pos_2nd_r  <= cfgdata_i[18:16];
      request_src_type_r <= cfgdata_i[21:20];
    end
  end

	//req_1(1)
	always @(posedge clk) begin
	  /* if(~rst_n) begin
	    request_addr_1st_row_r    <= 16'b0;
	    request_addr_1st_col_r    <= 14'b0;
	    request_addr_last_trans_r <= 1'b0;
	  end
	  else  */if(cfgreq_i && cfgfwd_i && (cfgid_i == 8'd1) && !cfgdata_i[31]) begin
	    request_addr_1st_row_r    <= cfgdata_i[15:0];
	    request_addr_1st_col_r    <= cfgdata_i[29:16];
	    request_addr_last_trans_r <= cfgdata_i[30];
	  end
	end
	
	//req_1(2)
	always @(posedge clk) begin
	  /* if(~rst_n)
	    request_cmd_access_addr_r   <= 20'b0;
	  else  */if(cfgreq_i && cfgfwd_i && (cfgid_i == 8'd1) && cfgdata_i[31])
	    request_cmd_access_addr_r   <= cfgdata_i[19:0];
	end
	
	/* �����жϵ�ǰ����������������ָ������ */
	always @(posedge clk) begin
	  /* if(~rst_n)
	    request_cmd_valid_r   <= 1'b0;
	  else  */if(cfgreq_i && cfgfwd_i && (cfgid_i == 8'd1) && cfgdata_i[31])
	    request_cmd_valid_r   <= 1'b1;
	  else if(request_valid_r)
	    request_cmd_valid_r   <= 1'b0;
	end
	
	
	
  //cfg info ----------------------------
  
  //cfg_0
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_ddr_channel_id_r <= 5'b0;
		cfg_VR_FR_r          <= 3'b0;
  		cfg_VR_id_r          <= 9'b0;
  		cfg_ch_cluster_num_r <= 3'b0;
  		cfg_D2D_flag_r       <= 1'b0;
  		cfg_read_write_r     <= 1'b0;
  		cfg_row_column_r     <= 1'b0;
  		cfg_broadcast_r      <= 1'b0;
  		cfg_stream_r         <= 1'b0;
      cfg_third_req_r      <= 1'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd0)) begin
  		cfg_ddr_channel_id_r <= cfgdata_i[ 4: 0];
		cfg_VR_FR_r          <= cfgdata_i[ 7: 5];
  		cfg_VR_id_r          <= cfgdata_i[16: 8];
  		cfg_ch_cluster_num_r <= cfgdata_i[22:20];
  		cfg_D2D_flag_r       <= cfgdata_i[26];
  		cfg_read_write_r     <= cfgdata_i[27];
  		cfg_row_column_r     <= cfgdata_i[28];
  		cfg_broadcast_r      <= cfgdata_i[29];
  		cfg_stream_r         <= cfgdata_i[30];
      cfg_third_req_r      <= cfgdata_i[31];
    end
  end
  
	
  //cfg_1
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_data_pos0_1st_r  <= 8'b0;
  		cfg_data_pos1_1st_r  <= 8'b0;
  		cfg_data_pos2_1st_r  <= 8'b0;
  		cfg_data_pos3_1st_r  <= 8'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd1)) begin
  		cfg_data_pos0_1st_r  <= cfgdata_i[ 7: 0];
  		cfg_data_pos1_1st_r  <= cfgdata_i[15: 8];
  		cfg_data_pos2_1st_r  <= cfgdata_i[23:16];
  		cfg_data_pos3_1st_r  <= cfgdata_i[31:24];
    end
  end
	
  //cfg_2
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_data_pos4_1st_r  <= 8'b0;
  		cfg_data_pos5_1st_r  <= 8'b0;
  		cfg_data_pos6_1st_r  <= 8'b0;
  		cfg_data_pos7_1st_r  <= 8'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd2)) begin
  		cfg_data_pos4_1st_r  <= cfgdata_i[ 7: 0];
  		cfg_data_pos5_1st_r  <= cfgdata_i[15: 8];
  		cfg_data_pos6_1st_r  <= cfgdata_i[23:16];
  		cfg_data_pos7_1st_r  <= cfgdata_i[31:24];
    end
  end
	
  //cfg_3
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_addr_pos0_1st_r  <= 8'b0;
  		cfg_addr_pos1_1st_r  <= 8'b0;
  		cfg_addr_pos2_1st_r  <= 8'b0;
  		cfg_addr_pos3_1st_r  <= 8'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd3)) begin
  		cfg_addr_pos0_1st_r  <= cfgdata_i[ 7: 0];
  		cfg_addr_pos1_1st_r  <= cfgdata_i[15: 8];
  		cfg_addr_pos2_1st_r  <= cfgdata_i[23:16];
  		cfg_addr_pos3_1st_r  <= cfgdata_i[31:24];
    end
  end
	
  //cfg_4
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_addr_pos4_1st_r  <= 8'b0;
  		cfg_addr_pos5_1st_r  <= 8'b0;
  		cfg_addr_pos6_1st_r  <= 8'b0;
  		cfg_addr_pos7_1st_r  <= 8'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd4)) begin
  		cfg_addr_pos4_1st_r  <= cfgdata_i[ 7: 0];
  		cfg_addr_pos5_1st_r  <= cfgdata_i[15: 8];
  		cfg_addr_pos6_1st_r  <= cfgdata_i[23:16];
  		cfg_addr_pos7_1st_r  <= cfgdata_i[31:24];
    end
  end
	
  //cfg_5
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_start_addr_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd5))
  		cfg_start_addr_r  <= cfgdata_i[29:0];
  end
	         //-----------------------------------------------------------// cfgid=5
             always@(posedge clk) begin                // cfgid=5
             	/* if(!rst_n) begin                                          // cfgid=5
             		pos_ok_start_pre_r <= 1'b0;                             // cfgid=5
               end                                                      // cfgid=5
               else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd5))      // cfgid=5
             		pos_ok_start_pre_r <= 1'b1;                             // cfgid=5
             	else                                                      // cfgid=5
             		pos_ok_start_pre_r <= 1'b0;                             // cfgid=5
             end                                                        // cfgid=5
	         //-----------------------------------------------------------// cfgid=5
	
  //cfg_6
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_row_num_1st_r    <= 16'b0;
  		cfg_column_num_1st_r <= 14'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd6)) begin
  		cfg_row_num_1st_r    <= cfgdata_i[15: 0];
  		cfg_column_num_1st_r <= cfgdata_i[29:16];
    end
  end
  
//	         //-----------------------------------------------------------// cfgid=6 
//             always@(posedge clk) begin                // cfgid=6 
//             	if(!rst_n) begin                                          // cfgid=6 
//             		pos_ok_start_en_r <= 1'b0;                              // cfgid=6 
//               end                                                      // cfgid=6 
//               else if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd6))      // cfgid=6 
//             		pos_ok_start_en_r <= 1'b1;                              // cfgid=6 
//             	else                                                      // cfgid=6 
//             		pos_ok_start_en_r <= 1'b0;                              // cfgid=6 
//             end                                                        // cfgid=6 
//	         //-----------------------------------------------------------// cfgid=6 
	
  //cfg_7
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_row_num_2nd_r    <= 16'b0;
  		cfg_column_num_2nd_r <= 14'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd7)) begin
  		cfg_row_num_2nd_r    <= cfgdata_i[15: 0];
  		cfg_column_num_2nd_r <= cfgdata_i[29:16];
    end
  end
	
  //cfg_8
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_data_pos0_2nd_r  <= 3'b0;
  		cfg_data_pos1_2nd_r  <= 3'b0;
  		cfg_data_pos2_2nd_r  <= 3'b0;
  		cfg_data_pos3_2nd_r  <= 3'b0;
  		cfg_data_pos4_2nd_r  <= 3'b0;
  		cfg_data_pos5_2nd_r  <= 3'b0;
  		cfg_data_pos6_2nd_r  <= 3'b0;
  		cfg_data_pos7_2nd_r  <= 3'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd8)) begin
  		cfg_data_pos0_2nd_r  <= cfgdata_i[ 2: 0];
  		cfg_data_pos1_2nd_r  <= cfgdata_i[ 5: 3];
  		cfg_data_pos2_2nd_r  <= cfgdata_i[ 8: 6];
  		cfg_data_pos3_2nd_r  <= cfgdata_i[11: 9];
  		cfg_data_pos4_2nd_r  <= cfgdata_i[14:12];
  		cfg_data_pos5_2nd_r  <= cfgdata_i[17:15];
  		cfg_data_pos6_2nd_r  <= cfgdata_i[20:18];
  		cfg_data_pos7_2nd_r  <= cfgdata_i[23:21];
    end
  end
	
  //cfg_9
  always@(posedge clk) begin
  	/* if(!rst_n) begin
  		cfg_addr_pos0_2nd_r  <= 3'b0;
  		cfg_addr_pos1_2nd_r  <= 3'b0;
  		cfg_addr_pos2_2nd_r  <= 3'b0;
  		cfg_addr_pos3_2nd_r  <= 3'b0;
  		cfg_addr_pos4_2nd_r  <= 3'b0;
  		cfg_addr_pos5_2nd_r  <= 3'b0;
  		cfg_addr_pos6_2nd_r  <= 3'b0;
  		cfg_addr_pos7_2nd_r  <= 3'b0;
    end
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd9)) begin
  		cfg_addr_pos0_2nd_r  <= cfgdata_i[ 2: 0];
  		cfg_addr_pos1_2nd_r  <= cfgdata_i[ 5: 3];
  		cfg_addr_pos2_2nd_r  <= cfgdata_i[ 8: 6];
  		cfg_addr_pos3_2nd_r  <= cfgdata_i[11: 9];
  		cfg_addr_pos4_2nd_r  <= cfgdata_i[14:12];
  		cfg_addr_pos5_2nd_r  <= cfgdata_i[17:15];
  		cfg_addr_pos6_2nd_r  <= cfgdata_i[20:18];
  		cfg_addr_pos7_2nd_r  <= cfgdata_i[23:21];
    end
  end
	
  //cfg_10
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_circu_times_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd10))
  		cfg_circu_times_r  <= cfgdata_i[29:0];
  end
	
  //cfg_11
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_col_addr_burst_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd11))
  		cfg_col_addr_burst_r  <= cfgdata_i[29:0];
  end
	
  //cfg_12
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_row_addr_burst_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd12))
  		cfg_row_addr_burst_r  <= cfgdata_i[29:0];
  end
	
  //cfg_13
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_2nd_addr_burst_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd13))
  		cfg_2nd_addr_burst_r  <= cfgdata_i[29:0];
  end
	
  //cfg_14
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_access_length_burst_r  <= 30'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd14))
  		cfg_access_length_burst_r  <= cfgdata_i[29:0];
  end
	
  //cfg_15
  always@(posedge clk) begin
  	/* if(!rst_n)
  		cfg_valid_r  <= 1'b0;
    else  */if(!cfgreq_i && cfgfwd_i && (cfgid_i == 8'd15))
  		cfg_valid_r  <= 1'b1;
  	else
  		cfg_valid_r  <= 1'b0;
  end
	
	
	
	//########################################
	// OUTPUT ---------- connection
	//########################################
	
  //request info
	assign	request_data_valid_o        = request_valid_r & !request_cmd_valid_r;
	assign	request_cmd_valid_o         = request_valid_r &  request_cmd_valid_r;
	assign	request_pos_1st_o           = request_pos_1st_r;
	assign	request_pos_2nd_o           = request_pos_2nd_r;
	assign	request_src_type_o          = request_src_type_r;
	assign	request_addr_1st_row_o      = request_addr_1st_row_r;
	assign	request_addr_1st_col_o      = request_addr_1st_col_r;
	assign	request_addr_last_trans_o   = request_addr_last_trans_r;
	assign	request_cmd_access_addr_o   = request_cmd_access_addr_r;
	//assign	request_mc_access_addr_o    = request_mc_access_addr_r;
	//assign	request_cop_access_addr_o   = request_mc_access_addr_r;
  

	//cfg info-------------------------------------------
	assign	cfg_valid_o           = cfg_valid_r;
//assign	cfg_get_clu_num_en_o  = cfg_get_clu_num_en_r;
//assign	cfg_pos_ok_en_o 			= cfg_pos_ok_en_r;
	
	assign	cfg_third_req_o       = cfg_third_req_r;
	assign	cfg_stream_o          = cfg_stream_r;
	assign	cfg_broadcast_o       = cfg_broadcast_r;
	assign	cfg_row_column_o      = cfg_row_column_r;
	assign	cfg_read_write_o      = cfg_read_write_r;
	assign	cfg_D2D_flag_o        = cfg_D2D_flag_r;
	assign	cfg_ch_cluster_num_o  = cfg_ch_cluster_num_r;
	assign	cfg_VR_id_o           = cfg_VR_id_r;
	assign  cfg_VR_FR_o           = cfg_VR_FR_r;
	assign	cfg_ddr_channel_id_o  = cfg_ddr_channel_id_r;
	
	
	//�����cfg info�����ߵ���ʽ�·���32��ddr_channel
	assign	cfg_data_pos0_1st_o  = cfg_data_pos0_1st_r;
	assign	cfg_data_pos1_1st_o  = cfg_data_pos1_1st_r;
	assign	cfg_data_pos2_1st_o  = cfg_data_pos2_1st_r;
	assign	cfg_data_pos3_1st_o  = cfg_data_pos3_1st_r;
	assign	cfg_data_pos4_1st_o  = cfg_data_pos4_1st_r;
	assign	cfg_data_pos5_1st_o  = cfg_data_pos5_1st_r;
	assign	cfg_data_pos6_1st_o  = cfg_data_pos6_1st_r;
	assign	cfg_data_pos7_1st_o  = cfg_data_pos7_1st_r;
	assign	cfg_data_pos0_2nd_o  = cfg_data_pos0_2nd_r;
	assign	cfg_data_pos1_2nd_o  = cfg_data_pos1_2nd_r;
	assign	cfg_data_pos2_2nd_o  = cfg_data_pos2_2nd_r;
	assign	cfg_data_pos3_2nd_o  = cfg_data_pos3_2nd_r;
	assign	cfg_data_pos4_2nd_o  = cfg_data_pos4_2nd_r;
	assign	cfg_data_pos5_2nd_o  = cfg_data_pos5_2nd_r;
	assign	cfg_data_pos6_2nd_o  = cfg_data_pos6_2nd_r;
	assign	cfg_data_pos7_2nd_o  = cfg_data_pos7_2nd_r;
	
	assign	cfg_addr_pos0_1st_o  = cfg_addr_pos0_1st_r;
	assign	cfg_addr_pos1_1st_o  = cfg_addr_pos1_1st_r;
	assign	cfg_addr_pos2_1st_o  = cfg_addr_pos2_1st_r;
	assign	cfg_addr_pos3_1st_o  = cfg_addr_pos3_1st_r;
	assign	cfg_addr_pos4_1st_o  = cfg_addr_pos4_1st_r;
	assign	cfg_addr_pos5_1st_o  = cfg_addr_pos5_1st_r;
	assign	cfg_addr_pos6_1st_o  = cfg_addr_pos6_1st_r;
	assign	cfg_addr_pos7_1st_o  = cfg_addr_pos7_1st_r;
	assign	cfg_addr_pos0_2nd_o  = cfg_addr_pos0_2nd_r;
	assign	cfg_addr_pos1_2nd_o  = cfg_addr_pos1_2nd_r;
	assign	cfg_addr_pos2_2nd_o  = cfg_addr_pos2_2nd_r;
	assign	cfg_addr_pos3_2nd_o  = cfg_addr_pos3_2nd_r;
	assign	cfg_addr_pos4_2nd_o  = cfg_addr_pos4_2nd_r;
	assign	cfg_addr_pos5_2nd_o  = cfg_addr_pos5_2nd_r;
	assign	cfg_addr_pos6_2nd_o  = cfg_addr_pos6_2nd_r;
	assign	cfg_addr_pos7_2nd_o  = cfg_addr_pos7_2nd_r;
	
	
	assign	cfg_start_addr_o     = cfg_start_addr_r;
	assign	cfg_row_num_1st_o    = cfg_row_num_1st_r;
	assign	cfg_column_num_1st_o = cfg_column_num_1st_r;
	assign	cfg_row_num_2nd_o    = cfg_row_num_2nd_r;
	assign	cfg_column_num_2nd_o = cfg_column_num_2nd_r;
	assign	cfg_circu_times_o    = cfg_circu_times_r;

	assign	cfg_col_addr_burst_o      = cfg_col_addr_burst_r;
	assign	cfg_row_addr_burst_o      = cfg_row_addr_burst_r;
	assign	cfg_2nd_addr_burst_o      = cfg_2nd_addr_burst_r;
	assign	cfg_access_length_burst_o = cfg_access_length_burst_r;
	
cfg_pos_ok_v2   cfg_pos_ok_v2(
    .clk(clk), 
  //  .rst_n(rst_n), 
    .cfg_broadcast_i      (cfg_broadcast_r), 
    .pos_ok_start_pre_i   (pos_ok_start_pre_r),    //����cfgid=5
   // .pos_ok_start_en_i    (pos_ok_start_en_r),     //����cfgid=6
    .cfg_row_column_i     (cfg_row_column_r),      //�������ȼ�   ����cfgid=0
    .cfg_ch_cluster_num_i (cfg_ch_cluster_num_r),  //���ôظ���   ����cfgid=0
    .cfg_row_num_1st_i    (cfg_row_num_1st_r),     //һ����������    ����cfgid=6
    .cfg_column_num_1st_i (cfg_column_num_1st_r),  //һ����������    ����cfgid=6
    
    .cfg_start_pos_row_0_o(cfg_start_pos_row_0_o), 
    .cfg_start_pos_col_0_o(cfg_start_pos_col_0_o), 
    .cfg_start_pos_row_1_o(cfg_start_pos_row_1_o), 
    .cfg_start_pos_col_1_o(cfg_start_pos_col_1_o), 
    .cfg_start_pos_row_2_o(cfg_start_pos_row_2_o), 
    .cfg_start_pos_col_2_o(cfg_start_pos_col_2_o), 
    .cfg_start_pos_row_3_o(cfg_start_pos_row_3_o), 
    .cfg_start_pos_col_3_o(cfg_start_pos_col_3_o), 
    .cfg_start_pos_row_4_o(cfg_start_pos_row_4_o), 
    .cfg_start_pos_col_4_o(cfg_start_pos_col_4_o), 
    .cfg_start_pos_row_5_o(cfg_start_pos_row_5_o), 
    .cfg_start_pos_col_5_o(cfg_start_pos_col_5_o), 
    .cfg_start_pos_row_6_o(cfg_start_pos_row_6_o), 
    .cfg_start_pos_col_6_o(cfg_start_pos_col_6_o), 
    .cfg_start_pos_row_7_o(cfg_start_pos_row_7_o), 
    .cfg_start_pos_col_7_o(cfg_start_pos_col_7_o)
    );
	
	

endmodule
