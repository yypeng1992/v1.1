interface my_if(input clk, input reset_n);

logic [7:0]data;
logic valid;

endinterface
